module main

fn main() {
	println('Hello from v lang!')
}
